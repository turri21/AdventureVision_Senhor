-------------------------------------------------------------------------------
--
-- The G port controller.
--
-- $Id: t400_io_g-c.vhd,v 1.1.1.1 2006/05/06 01:56:44 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_io_g_rtl_c0 of t400_io_g is

  for rtl
  end for;

end t400_io_g_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_io_g-c.vhd,v $
-- Revision 1.1.1.1  2006/05/06 01:56:44  arniml
-- import from local CVS repository, LOC_CVS_0_1
--
-------------------------------------------------------------------------------
