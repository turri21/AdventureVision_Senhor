-------------------------------------------------------------------------------
--
-- The timer unit.
--
-- $Id: t400_timer-c.vhd,v 1.1.1.1 2006/06/10 17:50:15 arnim Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_timer_rtl_c0 of t400_timer is

  for rtl
  end for;

end t400_timer_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_timer-c.vhd,v $
-- Revision 1.1.1.1  2006/06/10 17:50:15  arnim
-- copied from opencores.org repository, pre-1.0 release on 10-Jun-2006
--
-- Revision 1.1  2006/05/20 02:47:12  arniml
-- initial check-in
--
-------------------------------------------------------------------------------
