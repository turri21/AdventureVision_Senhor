-------------------------------------------------------------------------------
--
-- The stack unit.
--
-- $Id: t400_stack-c.vhd,v 1.1.1.1 2006/05/06 01:56:45 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_stack_rtl_c0 of t400_stack is

  for rtl
  end for;

end t400_stack_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_stack-c.vhd,v $
-- Revision 1.1.1.1  2006/05/06 01:56:45  arniml
-- import from local CVS repository, LOC_CVS_0_1
--
-------------------------------------------------------------------------------
