-------------------------------------------------------------------------------
--
-- The Arithmetic Logic Unit (ALU).
-- It contains the accumulator and the C flag.
--
-- $Id: t400_alu-c.vhd,v 1.1.1.1 2006/05/06 01:56:44 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_alu_rtl_c0 of t400_alu is

  for rtl
  end for;

end t400_alu_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_alu-c.vhd,v $
-- Revision 1.1.1.1  2006/05/06 01:56:44  arniml
-- import from local CVS repository, LOC_CVS_0_1
--
-------------------------------------------------------------------------------
