-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity adventurevision_bios is
	port(
		Clk	: in std_logic;
		A	: in std_logic_vector(9 downto 0);
		D	: out std_logic_vector(7 downto 0)
	);
end adventurevision_bios;

architecture rtl of adventurevision_bios is
	signal A_r : std_logic_vector(9 downto 0);
begin
	process (Clk)
	begin
		if Clk'event and Clk = '1' then
			A_r <= A;
		end if;
	end process;
	process (A_r)
	begin
		case to_integer(unsigned(A_r)) is
		when 000000 => D <= "11110101";	-- 0x0000
		when 000001 => D <= "00000100";	-- 0x0001
		when 000002 => D <= "00000000";	-- 0x0002
		when 000003 => D <= "00000100";	-- 0x0003
		when 000004 => D <= "00110110";	-- 0x0004
		when 000005 => D <= "00000100";	-- 0x0005
		when 000006 => D <= "01110001";	-- 0x0006
		when 000007 => D <= "00000100";	-- 0x0007
		when 000008 => D <= "11110000";	-- 0x0008
		when 000009 => D <= "00100100";	-- 0x0009
		when 000010 => D <= "10100000";	-- 0x000A
		when 000011 => D <= "01000100";	-- 0x000B
		when 000012 => D <= "10111001";	-- 0x000C
		when 000013 => D <= "01100100";	-- 0x000D
		when 000014 => D <= "01100001";	-- 0x000E
		when 000015 => D <= "01100100";	-- 0x000F
		when 000016 => D <= "00100100";	-- 0x0010
		when 000017 => D <= "01000100";	-- 0x0011
		when 000018 => D <= "11100010";	-- 0x0012
		when 000019 => D <= "01000100";	-- 0x0013
		when 000020 => D <= "11101111";	-- 0x0014
		when 000021 => D <= "00000100";	-- 0x0015
		when 000022 => D <= "00101011";	-- 0x0016
		when 000023 => D <= "01100100";	-- 0x0017
		when 000024 => D <= "10011010";	-- 0x0018
		when 000025 => D <= "01100100";	-- 0x0019
		when 000026 => D <= "11001110";	-- 0x001A
		when 000027 => D <= "01100100";	-- 0x001B
		when 000028 => D <= "10101001";	-- 0x001C
		when 000029 => D <= "01000100";	-- 0x001D
		when 000030 => D <= "11111111";	-- 0x001E
		when 000031 => D <= "01100100";	-- 0x001F
		when 000032 => D <= "00001110";	-- 0x0020
		when 000033 => D <= "01100100";	-- 0x0021
		when 000034 => D <= "00011101";	-- 0x0022
		when 000035 => D <= "00100100";	-- 0x0023
		when 000036 => D <= "10010111";	-- 0x0024
		when 000037 => D <= "01100100";	-- 0x0025
		when 000038 => D <= "11110001";	-- 0x0026
		when 000039 => D <= "01100100";	-- 0x0027
		when 000040 => D <= "11101111";	-- 0x0028
		when 000041 => D <= "01100100";	-- 0x0029
		when 000042 => D <= "11101101";	-- 0x002A
		when 000043 => D <= "10111000";	-- 0x002B
		when 000044 => D <= "00111111";	-- 0x002C
		when 000045 => D <= "10111001";	-- 0x002D
		when 000046 => D <= "00100000";	-- 0x002E
		when 000047 => D <= "00100111";	-- 0x002F
		when 000048 => D <= "10110000";	-- 0x0030
		when 000049 => D <= "00000000";	-- 0x0031
		when 000050 => D <= "11001000";	-- 0x0032
		when 000051 => D <= "11101001";	-- 0x0033
		when 000052 => D <= "00110000";	-- 0x0034
		when 000053 => D <= "10000011";	-- 0x0035
		when 000054 => D <= "11000101";	-- 0x0036
		when 000055 => D <= "10111000";	-- 0x0037
		when 000056 => D <= "00111111";	-- 0x0038
		when 000057 => D <= "00010000";	-- 0x0039
		when 000058 => D <= "01000110";	-- 0x003A
		when 000059 => D <= "00111010";	-- 0x003B
		when 000060 => D <= "01010110";	-- 0x003C
		when 000061 => D <= "00111100";	-- 0x003D
		when 000062 => D <= "10111001";	-- 0x003E
		when 000063 => D <= "00000001";	-- 0x003F
		when 000064 => D <= "11111001";	-- 0x0040
		when 000065 => D <= "00111001";	-- 0x0041
		when 000066 => D <= "10111000";	-- 0x0042
		when 000067 => D <= "00000101";	-- 0x0043
		when 000068 => D <= "00011000";	-- 0x0044
		when 000069 => D <= "11111000";	-- 0x0045
		when 000070 => D <= "10010110";	-- 0x0046
		when 000071 => D <= "01010000";	-- 0x0047
		when 000072 => D <= "00100111";	-- 0x0048
		when 000073 => D <= "00111010";	-- 0x0049
		when 000074 => D <= "00011001";	-- 0x004A
		when 000075 => D <= "11111001";	-- 0x004B
		when 000076 => D <= "01010010";	-- 0x004C
		when 000077 => D <= "01101101";	-- 0x004D
		when 000078 => D <= "00000100";	-- 0x004E
		when 000079 => D <= "01000001";	-- 0x004F
		when 000080 => D <= "00100011";	-- 0x0050
		when 000081 => D <= "00100000";	-- 0x0051
		when 000082 => D <= "00111010";	-- 0x0052
		when 000083 => D <= "10000000";	-- 0x0053
		when 000084 => D <= "00100011";	-- 0x0054
		when 000085 => D <= "01000000";	-- 0x0055
		when 000086 => D <= "00111010";	-- 0x0056
		when 000087 => D <= "00011000";	-- 0x0057
		when 000088 => D <= "10000000";	-- 0x0058
		when 000089 => D <= "00100011";	-- 0x0059
		when 000090 => D <= "01100000";	-- 0x005A
		when 000091 => D <= "00111010";	-- 0x005B
		when 000092 => D <= "00011000";	-- 0x005C
		when 000093 => D <= "10000000";	-- 0x005D
		when 000094 => D <= "00100011";	-- 0x005E
		when 000095 => D <= "10000000";	-- 0x005F
		when 000096 => D <= "00111010";	-- 0x0060
		when 000097 => D <= "00011000";	-- 0x0061
		when 000098 => D <= "10000000";	-- 0x0062
		when 000099 => D <= "00100011";	-- 0x0063
		when 000100 => D <= "10100000";	-- 0x0064
		when 000101 => D <= "00111010";	-- 0x0065
		when 000102 => D <= "00011000";	-- 0x0066
		when 000103 => D <= "10000000";	-- 0x0067
		when 000104 => D <= "00100011";	-- 0x0068
		when 000105 => D <= "00010000";	-- 0x0069
		when 000106 => D <= "00111010";	-- 0x006A
		when 000107 => D <= "00000100";	-- 0x006B
		when 000108 => D <= "01000100";	-- 0x006C
		when 000109 => D <= "00100111";	-- 0x006D
		when 000110 => D <= "00111001";	-- 0x006E
		when 000111 => D <= "11010101";	-- 0x006F
		when 000112 => D <= "10000011";	-- 0x0070
		when 000113 => D <= "00100111";	-- 0x0071
		when 000114 => D <= "00111001";	-- 0x0072
		when 000115 => D <= "11111001";	-- 0x0073
		when 000116 => D <= "01010011";	-- 0x0074
		when 000117 => D <= "11111000";	-- 0x0075
		when 000118 => D <= "00000011";	-- 0x0076
		when 000119 => D <= "00000011";	-- 0x0077
		when 000120 => D <= "10101001";	-- 0x0078
		when 000121 => D <= "10000001";	-- 0x0079
		when 000122 => D <= "00000011";	-- 0x007A
		when 000123 => D <= "11111100";	-- 0x007B
		when 000124 => D <= "11110110";	-- 0x007C
		when 000125 => D <= "10101001";	-- 0x007D
		when 000126 => D <= "11001001";	-- 0x007E
		when 000127 => D <= "11001001";	-- 0x007F
		when 000128 => D <= "10000001";	-- 0x0080
		when 000129 => D <= "10101010";	-- 0x0081
		when 000130 => D <= "11111001";	-- 0x0082
		when 000131 => D <= "11000101";	-- 0x0083
		when 000132 => D <= "10101000";	-- 0x0084
		when 000133 => D <= "00011000";	-- 0x0085
		when 000134 => D <= "10000000";	-- 0x0086
		when 000135 => D <= "10101001";	-- 0x0087
		when 000136 => D <= "00011000";	-- 0x0088
		when 000137 => D <= "10000000";	-- 0x0089
		when 000138 => D <= "10101010";	-- 0x008A
		when 000139 => D <= "00011000";	-- 0x008B
		when 000140 => D <= "10000000";	-- 0x008C
		when 000141 => D <= "10101011";	-- 0x008D
		when 000142 => D <= "11111011";	-- 0x008E
		when 000143 => D <= "00010111";	-- 0x008F
		when 000144 => D <= "10101110";	-- 0x0090
		when 000145 => D <= "11111010";	-- 0x0091
		when 000146 => D <= "10101101";	-- 0x0092
		when 000147 => D <= "10010110";	-- 0x0093
		when 000148 => D <= "10011111";	-- 0x0094
		when 000149 => D <= "10111110";	-- 0x0095
		when 000150 => D <= "00000110";	-- 0x0096
		when 000151 => D <= "00011101";	-- 0x0097
		when 000152 => D <= "11111101";	-- 0x0098
		when 000153 => D <= "00000011";	-- 0x0099
		when 000154 => D <= "11111100";	-- 0x009A
		when 000155 => D <= "10010110";	-- 0x009B
		when 000156 => D <= "10011111";	-- 0x009C
		when 000157 => D <= "10111101";	-- 0x009D
		when 000158 => D <= "00000001";	-- 0x009E
		when 000159 => D <= "10111111";	-- 0x009F
		when 000160 => D <= "00000000";	-- 0x00A0
		when 000161 => D <= "11110101";	-- 0x00A1
		when 000162 => D <= "00010100";	-- 0x00A2
		when 000163 => D <= "00000010";	-- 0x00A3
		when 000164 => D <= "11100101";	-- 0x00A4
		when 000165 => D <= "10101100";	-- 0x00A5
		when 000166 => D <= "00010111";	-- 0x00A6
		when 000167 => D <= "10010110";	-- 0x00A7
		when 000168 => D <= "10101101";	-- 0x00A8
		when 000169 => D <= "00100111";	-- 0x00A9
		when 000170 => D <= "00111001";	-- 0x00AA
		when 000171 => D <= "11010101";	-- 0x00AB
		when 000172 => D <= "10000011";	-- 0x00AC
		when 000173 => D <= "00110100";	-- 0x00AD
		when 000174 => D <= "01111000";	-- 0x00AE
		when 000175 => D <= "11111010";	-- 0x00AF
		when 000176 => D <= "00111001";	-- 0x00B0
		when 000177 => D <= "11111011";	-- 0x00B1
		when 000178 => D <= "10101000";	-- 0x00B2
		when 000179 => D <= "10000000";	-- 0x00B3
		when 000180 => D <= "00110111";	-- 0x00B4
		when 000181 => D <= "01011100";	-- 0x00B5
		when 000182 => D <= "11000110";	-- 0x00B6
		when 000183 => D <= "11000010";	-- 0x00B7
		when 000184 => D <= "00100011";	-- 0x00B8
		when 000185 => D <= "00000001";	-- 0x00B9
		when 000186 => D <= "10111000";	-- 0x00BA
		when 000187 => D <= "00111011";	-- 0x00BB
		when 000188 => D <= "01000000";	-- 0x00BC
		when 000189 => D <= "10100000";	-- 0x00BD
		when 000190 => D <= "00100111";	-- 0x00BE
		when 000191 => D <= "00111001";	-- 0x00BF
		when 000192 => D <= "00000100";	-- 0x00C0
		when 000193 => D <= "11001011";	-- 0x00C1
		when 000194 => D <= "11111101";	-- 0x00C2
		when 000195 => D <= "00111001";	-- 0x00C3
		when 000196 => D <= "11111110";	-- 0x00C4
		when 000197 => D <= "10101000";	-- 0x00C5
		when 000198 => D <= "10000000";	-- 0x00C6
		when 000199 => D <= "00110111";	-- 0x00C7
		when 000200 => D <= "01011111";	-- 0x00C8
		when 000201 => D <= "10010110";	-- 0x00C9
		when 000202 => D <= "10111000";	-- 0x00CA
		when 000203 => D <= "11111010";	-- 0x00CB
		when 000204 => D <= "00111001";	-- 0x00CC
		when 000205 => D <= "11111011";	-- 0x00CD
		when 000206 => D <= "10101000";	-- 0x00CE
		when 000207 => D <= "10000000";	-- 0x00CF
		when 000208 => D <= "00110111";	-- 0x00D0
		when 000209 => D <= "01001100";	-- 0x00D1
		when 000210 => D <= "00110111";	-- 0x00D2
		when 000211 => D <= "10010000";	-- 0x00D3
		when 000212 => D <= "11111101";	-- 0x00D4
		when 000213 => D <= "00111001";	-- 0x00D5
		when 000214 => D <= "11111110";	-- 0x00D6
		when 000215 => D <= "10101000";	-- 0x00D7
		when 000216 => D <= "10000000";	-- 0x00D8
		when 000217 => D <= "00110111";	-- 0x00D9
		when 000218 => D <= "01001111";	-- 0x00DA
		when 000219 => D <= "00110111";	-- 0x00DB
		when 000220 => D <= "10010000";	-- 0x00DC
		when 000221 => D <= "11111011";	-- 0x00DD
		when 000222 => D <= "00000011";	-- 0x00DE
		when 000223 => D <= "00000101";	-- 0x00DF
		when 000224 => D <= "10101011";	-- 0x00E0
		when 000225 => D <= "11100110";	-- 0x00E1
		when 000226 => D <= "11101110";	-- 0x00E2
		when 000227 => D <= "00000011";	-- 0x00E3
		when 000228 => D <= "00000110";	-- 0x00E4
		when 000229 => D <= "10101011";	-- 0x00E5
		when 000230 => D <= "00011010";	-- 0x00E6
		when 000231 => D <= "11111010";	-- 0x00E7
		when 000232 => D <= "00000011";	-- 0x00E8
		when 000233 => D <= "11111100";	-- 0x00E9
		when 000234 => D <= "10010110";	-- 0x00EA
		when 000235 => D <= "11101110";	-- 0x00EB
		when 000236 => D <= "10111010";	-- 0x00EC
		when 000237 => D <= "00000001";	-- 0x00ED
		when 000238 => D <= "00000100";	-- 0x00EE
		when 000239 => D <= "10001110";	-- 0x00EF
		when 000240 => D <= "00100111";	-- 0x00F0
		when 000241 => D <= "00111001";	-- 0x00F1
		when 000242 => D <= "11111001";	-- 0x00F2
		when 000243 => D <= "01010011";	-- 0x00F3
		when 000244 => D <= "11111000";	-- 0x00F4
		when 000245 => D <= "00000011";	-- 0x00F5
		when 000246 => D <= "00000011";	-- 0x00F6
		when 000247 => D <= "10101001";	-- 0x00F7
		when 000248 => D <= "10000001";	-- 0x00F8
		when 000249 => D <= "00000011";	-- 0x00F9
		when 000250 => D <= "11111100";	-- 0x00FA
		when 000251 => D <= "11100110";	-- 0x00FB
		when 000252 => D <= "11111111";	-- 0x00FC
		when 000253 => D <= "00100100";	-- 0x00FD
		when 000254 => D <= "00101011";	-- 0x00FE
		when 000255 => D <= "11001001";	-- 0x00FF
		when 000256 => D <= "11001001";	-- 0x0100
		when 000257 => D <= "10000001";	-- 0x0101
		when 000258 => D <= "10101010";	-- 0x0102
		when 000259 => D <= "11111001";	-- 0x0103
		when 000260 => D <= "11000101";	-- 0x0104
		when 000261 => D <= "10101000";	-- 0x0105
		when 000262 => D <= "00011000";	-- 0x0106
		when 000263 => D <= "10000000";	-- 0x0107
		when 000264 => D <= "10101001";	-- 0x0108
		when 000265 => D <= "00011000";	-- 0x0109
		when 000266 => D <= "10000000";	-- 0x010A
		when 000267 => D <= "10101010";	-- 0x010B
		when 000268 => D <= "00011000";	-- 0x010C
		when 000269 => D <= "10000000";	-- 0x010D
		when 000270 => D <= "10101011";	-- 0x010E
		when 000271 => D <= "11111011";	-- 0x010F
		when 000272 => D <= "00000011";	-- 0x0110
		when 000273 => D <= "00000001";	-- 0x0111
		when 000274 => D <= "10101110";	-- 0x0112
		when 000275 => D <= "11111010";	-- 0x0113
		when 000276 => D <= "10101101";	-- 0x0114
		when 000277 => D <= "11100110";	-- 0x0115
		when 000278 => D <= "00100001";	-- 0x0116
		when 000279 => D <= "10111110";	-- 0x0117
		when 000280 => D <= "00000110";	-- 0x0118
		when 000281 => D <= "00011101";	-- 0x0119
		when 000282 => D <= "11111101";	-- 0x011A
		when 000283 => D <= "00000011";	-- 0x011B
		when 000284 => D <= "11111100";	-- 0x011C
		when 000285 => D <= "10010110";	-- 0x011D
		when 000286 => D <= "00100001";	-- 0x011E
		when 000287 => D <= "10111101";	-- 0x011F
		when 000288 => D <= "00000001";	-- 0x0120
		when 000289 => D <= "10111111";	-- 0x0121
		when 000290 => D <= "00000000";	-- 0x0122
		when 000291 => D <= "11110101";	-- 0x0123
		when 000292 => D <= "00010100";	-- 0x0124
		when 000293 => D <= "00000010";	-- 0x0125
		when 000294 => D <= "11100101";	-- 0x0126
		when 000295 => D <= "10101100";	-- 0x0127
		when 000296 => D <= "00010111";	-- 0x0128
		when 000297 => D <= "10010110";	-- 0x0129
		when 000298 => D <= "00101111";	-- 0x012A
		when 000299 => D <= "00100111";	-- 0x012B
		when 000300 => D <= "00111001";	-- 0x012C
		when 000301 => D <= "11010101";	-- 0x012D
		when 000302 => D <= "10000011";	-- 0x012E
		when 000303 => D <= "00110100";	-- 0x012F
		when 000304 => D <= "01111000";	-- 0x0130
		when 000305 => D <= "10111000";	-- 0x0131
		when 000306 => D <= "00111000";	-- 0x0132
		when 000307 => D <= "11110000";	-- 0x0133
		when 000308 => D <= "01101011";	-- 0x0134
		when 000309 => D <= "10010110";	-- 0x0135
		when 000310 => D <= "01000001";	-- 0x0136
		when 000311 => D <= "00011000";	-- 0x0137
		when 000312 => D <= "11110000";	-- 0x0138
		when 000313 => D <= "01101010";	-- 0x0139
		when 000314 => D <= "10010110";	-- 0x013A
		when 000315 => D <= "01000001";	-- 0x013B
		when 000316 => D <= "00011000";	-- 0x013C
		when 000317 => D <= "11110000";	-- 0x013D
		when 000318 => D <= "01011100";	-- 0x013E
		when 000319 => D <= "10010110";	-- 0x013F
		when 000320 => D <= "01010001";	-- 0x0140
		when 000321 => D <= "10111000";	-- 0x0141
		when 000322 => D <= "00111000";	-- 0x0142
		when 000323 => D <= "11110000";	-- 0x0143
		when 000324 => D <= "01101110";	-- 0x0144
		when 000325 => D <= "10010110";	-- 0x0145
		when 000326 => D <= "01010111";	-- 0x0146
		when 000327 => D <= "00011000";	-- 0x0147
		when 000328 => D <= "11110000";	-- 0x0148
		when 000329 => D <= "01101101";	-- 0x0149
		when 000330 => D <= "10010110";	-- 0x014A
		when 000331 => D <= "01010111";	-- 0x014B
		when 000332 => D <= "00011000";	-- 0x014C
		when 000333 => D <= "11110000";	-- 0x014D
		when 000334 => D <= "01011111";	-- 0x014E
		when 000335 => D <= "11000110";	-- 0x014F
		when 000336 => D <= "01010111";	-- 0x0150
		when 000337 => D <= "00100011";	-- 0x0151
		when 000338 => D <= "00000010";	-- 0x0152
		when 000339 => D <= "10111000";	-- 0x0153
		when 000340 => D <= "00111011";	-- 0x0154
		when 000341 => D <= "01000000";	-- 0x0155
		when 000342 => D <= "10100000";	-- 0x0156
		when 000343 => D <= "11111010";	-- 0x0157
		when 000344 => D <= "00111001";	-- 0x0158
		when 000345 => D <= "11111011";	-- 0x0159
		when 000346 => D <= "10101000";	-- 0x015A
		when 000347 => D <= "10000000";	-- 0x015B
		when 000348 => D <= "01001100";	-- 0x015C
		when 000349 => D <= "10010000";	-- 0x015D
		when 000350 => D <= "11111101";	-- 0x015E
		when 000351 => D <= "00111001";	-- 0x015F
		when 000352 => D <= "11111110";	-- 0x0160
		when 000353 => D <= "10101000";	-- 0x0161
		when 000354 => D <= "10000000";	-- 0x0162
		when 000355 => D <= "01001111";	-- 0x0163
		when 000356 => D <= "10010000";	-- 0x0164
		when 000357 => D <= "11111011";	-- 0x0165
		when 000358 => D <= "00000011";	-- 0x0166
		when 000359 => D <= "00000101";	-- 0x0167
		when 000360 => D <= "10101011";	-- 0x0168
		when 000361 => D <= "11100110";	-- 0x0169
		when 000362 => D <= "00001111";	-- 0x016A
		when 000363 => D <= "00000011";	-- 0x016B
		when 000364 => D <= "00000110";	-- 0x016C
		when 000365 => D <= "10101011";	-- 0x016D
		when 000366 => D <= "00011010";	-- 0x016E
		when 000367 => D <= "11111010";	-- 0x016F
		when 000368 => D <= "00000011";	-- 0x0170
		when 000369 => D <= "11111100";	-- 0x0171
		when 000370 => D <= "10010110";	-- 0x0172
		when 000371 => D <= "01110110";	-- 0x0173
		when 000372 => D <= "10111010";	-- 0x0174
		when 000373 => D <= "00000001";	-- 0x0175
		when 000374 => D <= "00100100";	-- 0x0176
		when 000375 => D <= "00001111";	-- 0x0177
		when 000376 => D <= "11111001";	-- 0x0178
		when 000377 => D <= "10101000";	-- 0x0179
		when 000378 => D <= "11000110";	-- 0x017A
		when 000379 => D <= "10001001";	-- 0x017B
		when 000380 => D <= "00000011";	-- 0x017C
		when 000381 => D <= "11111100";	-- 0x017D
		when 000382 => D <= "11110110";	-- 0x017E
		when 000383 => D <= "10001010";	-- 0x017F
		when 000384 => D <= "10010111";	-- 0x0180
		when 000385 => D <= "11111100";	-- 0x0181
		when 000386 => D <= "11110111";	-- 0x0182
		when 000387 => D <= "10101100";	-- 0x0183
		when 000388 => D <= "11111111";	-- 0x0184
		when 000389 => D <= "11110111";	-- 0x0185
		when 000390 => D <= "10101111";	-- 0x0186
		when 000391 => D <= "11101000";	-- 0x0187
		when 000392 => D <= "10000000";	-- 0x0188
		when 000393 => D <= "10000011";	-- 0x0189
		when 000394 => D <= "00010111";	-- 0x018A
		when 000395 => D <= "10101000";	-- 0x018B
		when 000396 => D <= "11111100";	-- 0x018C
		when 000397 => D <= "01010011";	-- 0x018D
		when 000398 => D <= "00001111";	-- 0x018E
		when 000399 => D <= "01000111";	-- 0x018F
		when 000400 => D <= "00101100";	-- 0x0190
		when 000401 => D <= "01010011";	-- 0x0191
		when 000402 => D <= "11110000";	-- 0x0192
		when 000403 => D <= "01000111";	-- 0x0193
		when 000404 => D <= "10101111";	-- 0x0194
		when 000405 => D <= "00100100";	-- 0x0195
		when 000406 => D <= "10000111";	-- 0x0196
		when 000407 => D <= "10111001";	-- 0x0197
		when 000408 => D <= "11100001";	-- 0x0198
		when 000409 => D <= "11111000";	-- 0x0199
		when 000410 => D <= "10010001";	-- 0x019A
		when 000411 => D <= "01110100";	-- 0x019B
		when 000412 => D <= "00001110";	-- 0x019C
		when 000413 => D <= "00010100";	-- 0x019D
		when 000414 => D <= "01110001";	-- 0x019E
		when 000415 => D <= "10000011";	-- 0x019F
		when 000416 => D <= "11010101";	-- 0x01A0
		when 000417 => D <= "10111001";	-- 0x01A1
		when 000418 => D <= "00000000";	-- 0x01A2
		when 000419 => D <= "00100111";	-- 0x01A3
		when 000420 => D <= "00111001";	-- 0x01A4
		when 000421 => D <= "10000001";	-- 0x01A5
		when 000422 => D <= "10010110";	-- 0x01A6
		when 000423 => D <= "10110010";	-- 0x01A7
		when 000424 => D <= "11111001";	-- 0x01A8
		when 000425 => D <= "01010011";	-- 0x01A9
		when 000426 => D <= "11111000";	-- 0x01AA
		when 000427 => D <= "00000011";	-- 0x01AB
		when 000428 => D <= "00001000";	-- 0x01AC
		when 000429 => D <= "10101001";	-- 0x01AD
		when 000430 => D <= "10010110";	-- 0x01AE
		when 000431 => D <= "10100101";	-- 0x01AF
		when 000432 => D <= "01000100";	-- 0x01B0
		when 000433 => D <= "00011000";	-- 0x01B1
		when 000434 => D <= "11110101";	-- 0x01B2
		when 000435 => D <= "00010100";	-- 0x01B3
		when 000436 => D <= "00000110";	-- 0x01B4
		when 000437 => D <= "11100101";	-- 0x01B5
		when 000438 => D <= "11110010";	-- 0x01B6
		when 000439 => D <= "10101000";	-- 0x01B7
		when 000440 => D <= "10111000";	-- 0x01B8
		when 000441 => D <= "00111011";	-- 0x01B9
		when 000442 => D <= "10110000";	-- 0x01BA
		when 000443 => D <= "00000000";	-- 0x01BB
		when 000444 => D <= "00011001";	-- 0x01BC
		when 000445 => D <= "11110101";	-- 0x01BD
		when 000446 => D <= "00010100";	-- 0x01BE
		when 000447 => D <= "00001000";	-- 0x01BF
		when 000448 => D <= "11100101";	-- 0x01C0
		when 000449 => D <= "00010100";	-- 0x01C1
		when 000450 => D <= "11110000";	-- 0x01C2
		when 000451 => D <= "10111000";	-- 0x01C3
		when 000452 => D <= "00111011";	-- 0x01C4
		when 000453 => D <= "11110000";	-- 0x01C5
		when 000454 => D <= "10010110";	-- 0x01C6
		when 000455 => D <= "11010100";	-- 0x01C7
		when 000456 => D <= "11111001";	-- 0x01C8
		when 000457 => D <= "01010011";	-- 0x01C9
		when 000458 => D <= "11111000";	-- 0x01CA
		when 000459 => D <= "10101001";	-- 0x01CB
		when 000460 => D <= "10000001";	-- 0x01CC
		when 000461 => D <= "01010011";	-- 0x01CD
		when 000462 => D <= "00001111";	-- 0x01CE
		when 000463 => D <= "10101100";	-- 0x01CF
		when 000464 => D <= "01010100";	-- 0x01D0
		when 000465 => D <= "11111111";	-- 0x01D1
		when 000466 => D <= "00100100";	-- 0x01D2
		when 000467 => D <= "11100000";	-- 0x01D3
		when 000468 => D <= "10111000";	-- 0x01D4
		when 000469 => D <= "00111110";	-- 0x01D5
		when 000470 => D <= "11110000";	-- 0x01D6
		when 000471 => D <= "00010111";	-- 0x01D7
		when 000472 => D <= "10010110";	-- 0x01D8
		when 000473 => D <= "11001000";	-- 0x01D9
		when 000474 => D <= "11111001";	-- 0x01DA
		when 000475 => D <= "01010011";	-- 0x01DB
		when 000476 => D <= "11111000";	-- 0x01DC
		when 000477 => D <= "10100000";	-- 0x01DD
		when 000478 => D <= "00100100";	-- 0x01DE
		when 000479 => D <= "10101000";	-- 0x01DF
		when 000480 => D <= "10111010";	-- 0x01E0
		when 000481 => D <= "00000000";	-- 0x01E1
		when 000482 => D <= "10111011";	-- 0x01E2
		when 000483 => D <= "00000000";	-- 0x01E3
		when 000484 => D <= "01010100";	-- 0x01E4
		when 000485 => D <= "10111001";	-- 0x01E5
		when 000486 => D <= "11000110";	-- 0x01E6
		when 000487 => D <= "11101110";	-- 0x01E7
		when 000488 => D <= "11110101";	-- 0x01E8
		when 000489 => D <= "00010100";	-- 0x01E9
		when 000490 => D <= "00000100";	-- 0x01EA
		when 000491 => D <= "11100101";	-- 0x01EB
		when 000492 => D <= "00100100";	-- 0x01EC
		when 000493 => D <= "11100100";	-- 0x01ED
		when 000494 => D <= "11101100";	-- 0x01EE
		when 000495 => D <= "11100100";	-- 0x01EF
		when 000496 => D <= "11111010";	-- 0x01F0
		when 000497 => D <= "01110100";	-- 0x01F1
		when 000498 => D <= "01100001";	-- 0x01F2
		when 000499 => D <= "11111011";	-- 0x01F3
		when 000500 => D <= "01110100";	-- 0x01F4
		when 000501 => D <= "00100100";	-- 0x01F5
		when 000502 => D <= "11110101";	-- 0x01F6
		when 000503 => D <= "00010100";	-- 0x01F7
		when 000504 => D <= "00001010";	-- 0x01F8
		when 000505 => D <= "11100101";	-- 0x01F9
		when 000506 => D <= "01110100";	-- 0x01FA
		when 000507 => D <= "00001110";	-- 0x01FB
		when 000508 => D <= "11001001";	-- 0x01FC
		when 000509 => D <= "00010100";	-- 0x01FD
		when 000510 => D <= "01110001";	-- 0x01FE
		when 000511 => D <= "10111000";	-- 0x01FF
		when 000512 => D <= "00111011";	-- 0x0200
		when 000513 => D <= "11110000";	-- 0x0201
		when 000514 => D <= "10010110";	-- 0x0202
		when 000515 => D <= "00000110";	-- 0x0203
		when 000516 => D <= "00100100";	-- 0x0204
		when 000517 => D <= "10101000";	-- 0x0205
		when 000518 => D <= "10111000";	-- 0x0206
		when 000519 => D <= "00111100";	-- 0x0207
		when 000520 => D <= "11110000";	-- 0x0208
		when 000521 => D <= "01101001";	-- 0x0209
		when 000522 => D <= "11100110";	-- 0x020A
		when 000523 => D <= "00010110";	-- 0x020B
		when 000524 => D <= "10111000";	-- 0x020C
		when 000525 => D <= "00111110";	-- 0x020D
		when 000526 => D <= "11110000";	-- 0x020E
		when 000527 => D <= "00010111";	-- 0x020F
		when 000528 => D <= "10010110";	-- 0x0210
		when 000529 => D <= "00010110";	-- 0x0211
		when 000530 => D <= "11111001";	-- 0x0212
		when 000531 => D <= "01010011";	-- 0x0213
		when 000532 => D <= "11111000";	-- 0x0214
		when 000533 => D <= "10100000";	-- 0x0215
		when 000534 => D <= "00100100";	-- 0x0216
		when 000535 => D <= "10101000";	-- 0x0217
		when 000536 => D <= "10000001";	-- 0x0218
		when 000537 => D <= "10010110";	-- 0x0219
		when 000538 => D <= "00100100";	-- 0x021A
		when 000539 => D <= "11111001";	-- 0x021B
		when 000540 => D <= "01010011";	-- 0x021C
		when 000541 => D <= "11111000";	-- 0x021D
		when 000542 => D <= "00000011";	-- 0x021E
		when 000543 => D <= "00001000";	-- 0x021F
		when 000544 => D <= "10101001";	-- 0x0220
		when 000545 => D <= "10010110";	-- 0x0221
		when 000546 => D <= "00011000";	-- 0x0222
		when 000547 => D <= "10000011";	-- 0x0223
		when 000548 => D <= "11110010";	-- 0x0224
		when 000549 => D <= "00101000";	-- 0x0225
		when 000550 => D <= "01000100";	-- 0x0226
		when 000551 => D <= "00011011";	-- 0x0227
		when 000552 => D <= "01010011";	-- 0x0228
		when 000553 => D <= "00001111";	-- 0x0229
		when 000554 => D <= "10101100";	-- 0x022A
		when 000555 => D <= "01010100";	-- 0x022B
		when 000556 => D <= "11111111";	-- 0x022C
		when 000557 => D <= "11111101";	-- 0x022D
		when 000558 => D <= "10101000";	-- 0x022E
		when 000559 => D <= "00100011";	-- 0x022F
		when 000560 => D <= "00000001";	-- 0x0230
		when 000561 => D <= "11100111";	-- 0x0231
		when 000562 => D <= "11101000";	-- 0x0232
		when 000563 => D <= "00110001";	-- 0x0233
		when 000564 => D <= "10101010";	-- 0x0234
		when 000565 => D <= "11111110";	-- 0x0235
		when 000566 => D <= "00111001";	-- 0x0236
		when 000567 => D <= "11111111";	-- 0x0237
		when 000568 => D <= "10101000";	-- 0x0238
		when 000569 => D <= "10000000";	-- 0x0239
		when 000570 => D <= "01001010";	-- 0x023A
		when 000571 => D <= "10010000";	-- 0x023B
		when 000572 => D <= "00100111";	-- 0x023C
		when 000573 => D <= "00111001";	-- 0x023D
		when 000574 => D <= "10111010";	-- 0x023E
		when 000575 => D <= "00000000";	-- 0x023F
		when 000576 => D <= "10111011";	-- 0x0240
		when 000577 => D <= "00000000";	-- 0x0241
		when 000578 => D <= "01010100";	-- 0x0242
		when 000579 => D <= "10111001";	-- 0x0243
		when 000580 => D <= "11000110";	-- 0x0244
		when 000581 => D <= "01011100";	-- 0x0245
		when 000582 => D <= "00100011";	-- 0x0246
		when 000583 => D <= "11111000";	-- 0x0247
		when 000584 => D <= "01011001";	-- 0x0248
		when 000585 => D <= "00000011";	-- 0x0249
		when 000586 => D <= "00000001";	-- 0x024A
		when 000587 => D <= "10101001";	-- 0x024B
		when 000588 => D <= "10000001";	-- 0x024C
		when 000589 => D <= "00000111";	-- 0x024D
		when 000590 => D <= "10010001";	-- 0x024E
		when 000591 => D <= "11000110";	-- 0x024F
		when 000592 => D <= "01010111";	-- 0x0250
		when 000593 => D <= "11110101";	-- 0x0251
		when 000594 => D <= "00010100";	-- 0x0252
		when 000595 => D <= "00000100";	-- 0x0253
		when 000596 => D <= "11100101";	-- 0x0254
		when 000597 => D <= "01000100";	-- 0x0255
		when 000598 => D <= "01000010";	-- 0x0256
		when 000599 => D <= "11001001";	-- 0x0257
		when 000600 => D <= "00100111";	-- 0x0258
		when 000601 => D <= "10010001";	-- 0x0259
		when 000602 => D <= "01000100";	-- 0x025A
		when 000603 => D <= "00011011";	-- 0x025B
		when 000604 => D <= "11111010";	-- 0x025C
		when 000605 => D <= "01110100";	-- 0x025D
		when 000606 => D <= "01100001";	-- 0x025E
		when 000607 => D <= "11111011";	-- 0x025F
		when 000608 => D <= "01110100";	-- 0x0260
		when 000609 => D <= "00100100";	-- 0x0261
		when 000610 => D <= "11110101";	-- 0x0262
		when 000611 => D <= "00010100";	-- 0x0263
		when 000612 => D <= "00001100";	-- 0x0264
		when 000613 => D <= "11100101";	-- 0x0265
		when 000614 => D <= "11111101";	-- 0x0266
		when 000615 => D <= "00010111";	-- 0x0267
		when 000616 => D <= "10101010";	-- 0x0268
		when 000617 => D <= "00100011";	-- 0x0269
		when 000618 => D <= "00000001";	-- 0x026A
		when 000619 => D <= "01000100";	-- 0x026B
		when 000620 => D <= "01101110";	-- 0x026C
		when 000621 => D <= "11100111";	-- 0x026D
		when 000622 => D <= "11101010";	-- 0x026E
		when 000623 => D <= "01101101";	-- 0x026F
		when 000624 => D <= "10101010";	-- 0x0270
		when 000625 => D <= "11111111";	-- 0x0271
		when 000626 => D <= "10101000";	-- 0x0272
		when 000627 => D <= "11111110";	-- 0x0273
		when 000628 => D <= "00111001";	-- 0x0274
		when 000629 => D <= "10000000";	-- 0x0275
		when 000630 => D <= "10101011";	-- 0x0276
		when 000631 => D <= "01001010";	-- 0x0277
		when 000632 => D <= "10010000";	-- 0x0278
		when 000633 => D <= "11111011";	-- 0x0279
		when 000634 => D <= "00110111";	-- 0x027A
		when 000635 => D <= "01011010";	-- 0x027B
		when 000636 => D <= "10010110";	-- 0x027C
		when 000637 => D <= "10001100";	-- 0x027D
		when 000638 => D <= "11101100";	-- 0x027E
		when 000639 => D <= "00111100";	-- 0x027F
		when 000640 => D <= "11111010";	-- 0x0280
		when 000641 => D <= "10000000";	-- 0x0281
		when 000642 => D <= "00110111";	-- 0x0282
		when 000643 => D <= "01001010";	-- 0x0283
		when 000644 => D <= "00110111";	-- 0x0284
		when 000645 => D <= "10010000";	-- 0x0285
		when 000646 => D <= "00100111";	-- 0x0286
		when 000647 => D <= "00111001";	-- 0x0287
		when 000648 => D <= "01110100";	-- 0x0288
		when 000649 => D <= "00001110";	-- 0x0289
		when 000650 => D <= "01000100";	-- 0x028A
		when 000651 => D <= "00011011";	-- 0x028B
		when 000652 => D <= "00100111";	-- 0x028C
		when 000653 => D <= "00111001";	-- 0x028D
		when 000654 => D <= "00100011";	-- 0x028E
		when 000655 => D <= "11111000";	-- 0x028F
		when 000656 => D <= "01011001";	-- 0x0290
		when 000657 => D <= "10101001";	-- 0x0291
		when 000658 => D <= "10000001";	-- 0x0292
		when 000659 => D <= "10101011";	-- 0x0293
		when 000660 => D <= "11111110";	-- 0x0294
		when 000661 => D <= "00111001";	-- 0x0295
		when 000662 => D <= "11111011";	-- 0x0296
		when 000663 => D <= "01010011";	-- 0x0297
		when 000664 => D <= "00110000";	-- 0x0298
		when 000665 => D <= "11000110";	-- 0x0299
		when 000666 => D <= "01111110";	-- 0x029A
		when 000667 => D <= "00101000";	-- 0x029B
		when 000668 => D <= "10101011";	-- 0x029C
		when 000669 => D <= "11111000";	-- 0x029D
		when 000670 => D <= "10111000";	-- 0x029E
		when 000671 => D <= "00110111";	-- 0x029F
		when 000672 => D <= "10100000";	-- 0x02A0
		when 000673 => D <= "00011000";	-- 0x02A1
		when 000674 => D <= "11111111";	-- 0x02A2
		when 000675 => D <= "00110111";	-- 0x02A3
		when 000676 => D <= "00010111";	-- 0x02A4
		when 000677 => D <= "10100000";	-- 0x02A5
		when 000678 => D <= "00011000";	-- 0x02A6
		when 000679 => D <= "11111110";	-- 0x02A7
		when 000680 => D <= "00110111";	-- 0x02A8
		when 000681 => D <= "00010111";	-- 0x02A9
		when 000682 => D <= "10100000";	-- 0x02AA
		when 000683 => D <= "11111101";	-- 0x02AB
		when 000684 => D <= "10101000";	-- 0x02AC
		when 000685 => D <= "00100011";	-- 0x02AD
		when 000686 => D <= "00000001";	-- 0x02AE
		when 000687 => D <= "11100111";	-- 0x02AF
		when 000688 => D <= "11101000";	-- 0x02B0
		when 000689 => D <= "10101111";	-- 0x02B1
		when 000690 => D <= "10111000";	-- 0x02B2
		when 000691 => D <= "00111010";	-- 0x02B3
		when 000692 => D <= "10100000";	-- 0x02B4
		when 000693 => D <= "11111011";	-- 0x02B5
		when 000694 => D <= "10101000";	-- 0x02B6
		when 000695 => D <= "01000100";	-- 0x02B7
		when 000696 => D <= "01111110";	-- 0x02B8
		when 000697 => D <= "00100011";	-- 0x02B9
		when 000698 => D <= "11111000";	-- 0x02BA
		when 000699 => D <= "01011001";	-- 0x02BB
		when 000700 => D <= "00000011";	-- 0x02BC
		when 000701 => D <= "00000101";	-- 0x02BD
		when 000702 => D <= "10101001";	-- 0x02BE
		when 000703 => D <= "10000001";	-- 0x02BF
		when 000704 => D <= "11000110";	-- 0x02C0
		when 000705 => D <= "11011011";	-- 0x02C1
		when 000706 => D <= "11110010";	-- 0x02C2
		when 000707 => D <= "11001000";	-- 0x02C3
		when 000708 => D <= "00011010";	-- 0x02C4
		when 000709 => D <= "00000111";	-- 0x02C5
		when 000710 => D <= "01000100";	-- 0x02C6
		when 000711 => D <= "11001010";	-- 0x02C7
		when 000712 => D <= "11001010";	-- 0x02C8
		when 000713 => D <= "00010111";	-- 0x02C9
		when 000714 => D <= "10010001";	-- 0x02CA
		when 000715 => D <= "00011001";	-- 0x02CB
		when 000716 => D <= "10000001";	-- 0x02CC
		when 000717 => D <= "10010110";	-- 0x02CD
		when 000718 => D <= "11010000";	-- 0x02CE
		when 000719 => D <= "10000011";	-- 0x02CF
		when 000720 => D <= "11110010";	-- 0x02D0
		when 000721 => D <= "11010110";	-- 0x02D1
		when 000722 => D <= "00011011";	-- 0x02D2
		when 000723 => D <= "00000111";	-- 0x02D3
		when 000724 => D <= "01000100";	-- 0x02D4
		when 000725 => D <= "11011000";	-- 0x02D5
		when 000726 => D <= "11001011";	-- 0x02D6
		when 000727 => D <= "00010111";	-- 0x02D7
		when 000728 => D <= "10010001";	-- 0x02D8
		when 000729 => D <= "00100111";	-- 0x02D9
		when 000730 => D <= "10000011";	-- 0x02DA
		when 000731 => D <= "00011001";	-- 0x02DB
		when 000732 => D <= "10000001";	-- 0x02DC
		when 000733 => D <= "10010110";	-- 0x02DD
		when 000734 => D <= "11010000";	-- 0x02DE
		when 000735 => D <= "00100011";	-- 0x02DF
		when 000736 => D <= "11111111";	-- 0x02E0
		when 000737 => D <= "10000011";	-- 0x02E1
		when 000738 => D <= "10111000";	-- 0x02E2
		when 000739 => D <= "00000000";	-- 0x02E3
		when 000740 => D <= "10111011";	-- 0x02E4
		when 000741 => D <= "00000100";	-- 0x02E5
		when 000742 => D <= "11111011";	-- 0x02E6
		when 000743 => D <= "00000111";	-- 0x02E7
		when 000744 => D <= "00111001";	-- 0x02E8
		when 000745 => D <= "00100111";	-- 0x02E9
		when 000746 => D <= "10010000";	-- 0x02EA
		when 000747 => D <= "11101000";	-- 0x02EB
		when 000748 => D <= "11101010";	-- 0x02EC
		when 000749 => D <= "11101011";	-- 0x02ED
		when 000750 => D <= "11100110";	-- 0x02EE
		when 000751 => D <= "10111000";	-- 0x02EF
		when 000752 => D <= "00000000";	-- 0x02F0
		when 000753 => D <= "10111011";	-- 0x02F1
		when 000754 => D <= "00000011";	-- 0x02F2
		when 000755 => D <= "11111011";	-- 0x02F3
		when 000756 => D <= "00111001";	-- 0x02F4
		when 000757 => D <= "00100011";	-- 0x02F5
		when 000758 => D <= "11111111";	-- 0x02F6
		when 000759 => D <= "10010000";	-- 0x02F7
		when 000760 => D <= "11101000";	-- 0x02F8
		when 000761 => D <= "11110111";	-- 0x02F9
		when 000762 => D <= "11101011";	-- 0x02FA
		when 000763 => D <= "11110011";	-- 0x02FB
		when 000764 => D <= "00100111";	-- 0x02FC
		when 000765 => D <= "00111001";	-- 0x02FD
		when 000766 => D <= "10000011";	-- 0x02FE
		when 000767 => D <= "11111001";	-- 0x02FF
		when 000768 => D <= "01010011";	-- 0x0300
		when 000769 => D <= "11111000";	-- 0x0301
		when 000770 => D <= "00000011";	-- 0x0302
		when 000771 => D <= "00000010";	-- 0x0303
		when 000772 => D <= "10101001";	-- 0x0304
		when 000773 => D <= "10000001";	-- 0x0305
		when 000774 => D <= "10101101";	-- 0x0306
		when 000775 => D <= "00011001";	-- 0x0307
		when 000776 => D <= "10000001";	-- 0x0308
		when 000777 => D <= "10101110";	-- 0x0309
		when 000778 => D <= "00011001";	-- 0x030A
		when 000779 => D <= "10000001";	-- 0x030B
		when 000780 => D <= "10101111";	-- 0x030C
		when 000781 => D <= "10000011";	-- 0x030D
		when 000782 => D <= "11111001";	-- 0x030E
		when 000783 => D <= "01010011";	-- 0x030F
		when 000784 => D <= "11111000";	-- 0x0310
		when 000785 => D <= "00000011";	-- 0x0311
		when 000786 => D <= "00000010";	-- 0x0312
		when 000787 => D <= "10101001";	-- 0x0313
		when 000788 => D <= "11111101";	-- 0x0314
		when 000789 => D <= "10010001";	-- 0x0315
		when 000790 => D <= "00011001";	-- 0x0316
		when 000791 => D <= "11111110";	-- 0x0317
		when 000792 => D <= "10010001";	-- 0x0318
		when 000793 => D <= "00011001";	-- 0x0319
		when 000794 => D <= "11111111";	-- 0x031A
		when 000795 => D <= "10010001";	-- 0x031B
		when 000796 => D <= "10000011";	-- 0x031C
		when 000797 => D <= "01110100";	-- 0x031D
		when 000798 => D <= "00001110";	-- 0x031E
		when 000799 => D <= "00100111";	-- 0x031F
		when 000800 => D <= "10010001";	-- 0x0320
		when 000801 => D <= "00011001";	-- 0x0321
		when 000802 => D <= "10010001";	-- 0x0322
		when 000803 => D <= "10000011";	-- 0x0323
		when 000804 => D <= "10111000";	-- 0x0324
		when 000805 => D <= "00101110";	-- 0x0325
		when 000806 => D <= "01101101";	-- 0x0326
		when 000807 => D <= "10101101";	-- 0x0327
		when 000808 => D <= "11110010";	-- 0x0328
		when 000809 => D <= "01001100";	-- 0x0329
		when 000810 => D <= "01010011";	-- 0x032A
		when 000811 => D <= "11111000";	-- 0x032B
		when 000812 => D <= "10010110";	-- 0x032C
		when 000813 => D <= "00101111";	-- 0x032D
		when 000814 => D <= "10000011";	-- 0x032E
		when 000815 => D <= "11111101";	-- 0x032F
		when 000816 => D <= "00000011";	-- 0x0330
		when 000817 => D <= "11111000";	-- 0x0331
		when 000818 => D <= "10101101";	-- 0x0332
		when 000819 => D <= "00011111";	-- 0x0333
		when 000820 => D <= "11111111";	-- 0x0334
		when 000821 => D <= "10010110";	-- 0x0335
		when 000822 => D <= "01000000";	-- 0x0336
		when 000823 => D <= "10111111";	-- 0x0337
		when 000824 => D <= "00000110";	-- 0x0338
		when 000825 => D <= "00011110";	-- 0x0339
		when 000826 => D <= "11111110";	-- 0x033A
		when 000827 => D <= "00110111";	-- 0x033B
		when 000828 => D <= "00010111";	-- 0x033C
		when 000829 => D <= "01100000";	-- 0x033D
		when 000830 => D <= "11100110";	-- 0x033E
		when 000831 => D <= "01000011";	-- 0x033F
		when 000832 => D <= "11111101";	-- 0x0340
		when 000833 => D <= "01100100";	-- 0x0341
		when 000834 => D <= "00101010";	-- 0x0342
		when 000835 => D <= "10111110";	-- 0x0343
		when 000836 => D <= "00000001";	-- 0x0344
		when 000837 => D <= "01100100";	-- 0x0345
		when 000838 => D <= "01000000";	-- 0x0346
		when 000839 => D <= "01010011";	-- 0x0347
		when 000840 => D <= "11111000";	-- 0x0348
		when 000841 => D <= "10010110";	-- 0x0349
		when 000842 => D <= "01001100";	-- 0x034A
		when 000843 => D <= "10000011";	-- 0x034B
		when 000844 => D <= "11111101";	-- 0x034C
		when 000845 => D <= "00000011";	-- 0x034D
		when 000846 => D <= "00001000";	-- 0x034E
		when 000847 => D <= "10101101";	-- 0x034F
		when 000848 => D <= "11001111";	-- 0x0350
		when 000849 => D <= "11111111";	-- 0x0351
		when 000850 => D <= "00000011";	-- 0x0352
		when 000851 => D <= "11111010";	-- 0x0353
		when 000852 => D <= "11100110";	-- 0x0354
		when 000853 => D <= "01011001";	-- 0x0355
		when 000854 => D <= "11111101";	-- 0x0356
		when 000855 => D <= "01100100";	-- 0x0357
		when 000856 => D <= "01000111";	-- 0x0358
		when 000857 => D <= "10111111";	-- 0x0359
		when 000858 => D <= "11111111";	-- 0x035A
		when 000859 => D <= "11101110";	-- 0x035B
		when 000860 => D <= "01010110";	-- 0x035C
		when 000861 => D <= "11110000";	-- 0x035D
		when 000862 => D <= "10101110";	-- 0x035E
		when 000863 => D <= "01100100";	-- 0x035F
		when 000864 => D <= "01010110";	-- 0x0360
		when 000865 => D <= "11110010";	-- 0x0361
		when 000866 => D <= "10000101";	-- 0x0362
		when 000867 => D <= "10101000";	-- 0x0363
		when 000868 => D <= "11100111";	-- 0x0364
		when 000869 => D <= "11100111";	-- 0x0365
		when 000870 => D <= "01101000";	-- 0x0366
		when 000871 => D <= "10101000";	-- 0x0367
		when 000872 => D <= "01101111";	-- 0x0368
		when 000873 => D <= "10101111";	-- 0x0369
		when 000874 => D <= "11110110";	-- 0x036A
		when 000875 => D <= "01110101";	-- 0x036B
		when 000876 => D <= "10000011";	-- 0x036C
		when 000877 => D <= "10101111";	-- 0x036D
		when 000878 => D <= "11101110";	-- 0x036E
		when 000879 => D <= "01110100";	-- 0x036F
		when 000880 => D <= "10111000";	-- 0x0370
		when 000881 => D <= "00101110";	-- 0x0371
		when 000882 => D <= "11110000";	-- 0x0372
		when 000883 => D <= "10101110";	-- 0x0373
		when 000884 => D <= "10000011";	-- 0x0374
		when 000885 => D <= "00000011";	-- 0x0375
		when 000886 => D <= "00000110";	-- 0x0376
		when 000887 => D <= "10101111";	-- 0x0377
		when 000888 => D <= "00011110";	-- 0x0378
		when 000889 => D <= "11111110";	-- 0x0379
		when 000890 => D <= "10111000";	-- 0x037A
		when 000891 => D <= "00101110";	-- 0x037B
		when 000892 => D <= "00110111";	-- 0x037C
		when 000893 => D <= "00010111";	-- 0x037D
		when 000894 => D <= "01100000";	-- 0x037E
		when 000895 => D <= "11100110";	-- 0x037F
		when 000896 => D <= "10000010";	-- 0x0380
		when 000897 => D <= "10000011";	-- 0x0381
		when 000898 => D <= "10111110";	-- 0x0382
		when 000899 => D <= "00000001";	-- 0x0383
		when 000900 => D <= "10000011";	-- 0x0384
		when 000901 => D <= "00110111";	-- 0x0385
		when 000902 => D <= "00010111";	-- 0x0386
		when 000903 => D <= "10101000";	-- 0x0387
		when 000904 => D <= "11100111";	-- 0x0388
		when 000905 => D <= "11100111";	-- 0x0389
		when 000906 => D <= "01101000";	-- 0x038A
		when 000907 => D <= "00110111";	-- 0x038B
		when 000908 => D <= "00010111";	-- 0x038C
		when 000909 => D <= "01101111";	-- 0x038D
		when 000910 => D <= "11100110";	-- 0x038E
		when 000911 => D <= "10010110";	-- 0x038F
		when 000912 => D <= "10101111";	-- 0x0390
		when 000913 => D <= "00000011";	-- 0x0391
		when 000914 => D <= "11111010";	-- 0x0392
		when 000915 => D <= "11100110";	-- 0x0393
		when 000916 => D <= "01101101";	-- 0x0394
		when 000917 => D <= "10000011";	-- 0x0395
		when 000918 => D <= "00000011";	-- 0x0396
		when 000919 => D <= "11111010";	-- 0x0397
		when 000920 => D <= "01100100";	-- 0x0398
		when 000921 => D <= "01101101";	-- 0x0399
		when 000922 => D <= "10111000";	-- 0x039A
		when 000923 => D <= "00110100";	-- 0x039B
		when 000924 => D <= "01100000";	-- 0x039C
		when 000925 => D <= "01010111";	-- 0x039D
		when 000926 => D <= "10100000";	-- 0x039E
		when 000927 => D <= "11110110";	-- 0x039F
		when 000928 => D <= "10100010";	-- 0x03A0
		when 000929 => D <= "10000011";	-- 0x03A1
		when 000930 => D <= "11001000";	-- 0x03A2
		when 000931 => D <= "11110000";	-- 0x03A3
		when 000932 => D <= "00000011";	-- 0x03A4
		when 000933 => D <= "00000001";	-- 0x03A5
		when 000934 => D <= "01010111";	-- 0x03A6
		when 000935 => D <= "10100000";	-- 0x03A7
		when 000936 => D <= "10000011";	-- 0x03A8
		when 000937 => D <= "00100011";	-- 0x03A9
		when 000938 => D <= "11000000";	-- 0x03AA
		when 000939 => D <= "00111010";	-- 0x03AB
		when 000940 => D <= "00100011";	-- 0x03AC
		when 000941 => D <= "00000001";	-- 0x03AD
		when 000942 => D <= "00111001";	-- 0x03AE
		when 000943 => D <= "10111000";	-- 0x03AF
		when 000944 => D <= "00000000";	-- 0x03B0
		when 000945 => D <= "00100111";	-- 0x03B1
		when 000946 => D <= "10010000";	-- 0x03B2
		when 000947 => D <= "10000000";	-- 0x03B3
		when 000948 => D <= "10111010";	-- 0x03B4
		when 000949 => D <= "00010100";	-- 0x03B5
		when 000950 => D <= "11101010";	-- 0x03B6
		when 000951 => D <= "10110110";	-- 0x03B7
		when 000952 => D <= "00000000";	-- 0x03B8
		when 000953 => D <= "00100011";	-- 0x03B9
		when 000954 => D <= "00000001";	-- 0x03BA
		when 000955 => D <= "10010000";	-- 0x03BB
		when 000956 => D <= "10000000";	-- 0x03BC
		when 000957 => D <= "11111001";	-- 0x03BD
		when 000958 => D <= "00111010";	-- 0x03BE
		when 000959 => D <= "10111010";	-- 0x03BF
		when 000960 => D <= "00100110";	-- 0x03C0
		when 000961 => D <= "11101010";	-- 0x03C1
		when 000962 => D <= "11000001";	-- 0x03C2
		when 000963 => D <= "00000000";	-- 0x03C3
		when 000964 => D <= "01000111";	-- 0x03C4
		when 000965 => D <= "00111010";	-- 0x03C5
		when 000966 => D <= "10111010";	-- 0x03C6
		when 000967 => D <= "00100001";	-- 0x03C7
		when 000968 => D <= "11101010";	-- 0x03C8
		when 000969 => D <= "11001000";	-- 0x03C9
		when 000970 => D <= "00100111";	-- 0x03CA
		when 000971 => D <= "00111001";	-- 0x03CB
		when 000972 => D <= "00111010";	-- 0x03CC
		when 000973 => D <= "10000011";	-- 0x03CD
		when 000974 => D <= "00100111";	-- 0x03CE
		when 000975 => D <= "00111001";	-- 0x03CF
		when 000976 => D <= "10111000";	-- 0x03D0
		when 000977 => D <= "00000001";	-- 0x03D1
		when 000978 => D <= "00100111";	-- 0x03D2
		when 000979 => D <= "10010000";	-- 0x03D3
		when 000980 => D <= "11111101";	-- 0x03D4
		when 000981 => D <= "00011000";	-- 0x03D5
		when 000982 => D <= "10010000";	-- 0x03D6
		when 000983 => D <= "11111110";	-- 0x03D7
		when 000984 => D <= "00011000";	-- 0x03D8
		when 000985 => D <= "10010000";	-- 0x03D9
		when 000986 => D <= "11111111";	-- 0x03DA
		when 000987 => D <= "00011000";	-- 0x03DB
		when 000988 => D <= "10010000";	-- 0x03DC
		when 000989 => D <= "11010101";	-- 0x03DD
		when 000990 => D <= "10111001";	-- 0x03DE
		when 000991 => D <= "00000001";	-- 0x03DF
		when 000992 => D <= "00010100";	-- 0x03E0
		when 000993 => D <= "01110001";	-- 0x03E1
		when 000994 => D <= "00010100";	-- 0x03E2
		when 000995 => D <= "00110110";	-- 0x03E3
		when 000996 => D <= "00100011";	-- 0x03E4
		when 000997 => D <= "11111000";	-- 0x03E5
		when 000998 => D <= "00111001";	-- 0x03E6
		when 000999 => D <= "00001001";	-- 0x03E7
		when 001000 => D <= "01110010";	-- 0x03E8
		when 001001 => D <= "11100010";	-- 0x03E9
		when 001002 => D <= "11110101";	-- 0x03EA
		when 001003 => D <= "00000100";	-- 0x03EB
		when 001004 => D <= "00000000";	-- 0x03EC
		when 001005 => D <= "00111100";	-- 0x03ED
		when 001006 => D <= "10000011";	-- 0x03EE
		when 001007 => D <= "00111101";	-- 0x03EF
		when 001008 => D <= "10000011";	-- 0x03F0
		when 001009 => D <= "11111101";	-- 0x03F1
		when 001010 => D <= "00010111";	-- 0x03F2
		when 001011 => D <= "10101001";	-- 0x03F3
		when 001012 => D <= "00100011";	-- 0x03F4
		when 001013 => D <= "10000000";	-- 0x03F5
		when 001014 => D <= "11100111";	-- 0x03F6
		when 001015 => D <= "11101001";	-- 0x03F7
		when 001016 => D <= "11110110";	-- 0x03F8
		when 001017 => D <= "10000011";	-- 0x03F9
		when 001018 => D <= "00110000";	-- 0x03FA
		when 001019 => D <= "00101001";	-- 0x03FB
		when 001020 => D <= "01011100";	-- 0x03FC
		when 001021 => D <= "00110010";	-- 0x03FD
		when 001022 => D <= "00110101";	-- 0x03FE
		when 001023 => D <= "00110110";	-- 0x03FF
		when others => D <= "--------";
		end case;
	end process;
end;
