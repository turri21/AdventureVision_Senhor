-------------------------------------------------------------------------------
--
-- The IN port controller.
--
-- $Id: t400_io_in-c.vhd,v 1.1.1.1 2006/06/10 17:50:15 arnim Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_io_in_rtl_c0 of t400_io_in is

  for rtl
  end for;

end t400_io_in_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_io_in-c.vhd,v $
-- Revision 1.1.1.1  2006/06/10 17:50:15  arnim
-- copied from opencores.org repository, pre-1.0 release on 10-Jun-2006
--
-- Revision 1.1  2006/05/22 00:00:55  arniml
-- initial check-in
--
-------------------------------------------------------------------------------
