-------------------------------------------------------------------------------
--
-- The clock generation unit.
-- PHI1 clock and input/output clock enables are generated here.
--
-- $Id: t400_clkgen-c.vhd,v 1.1.1.1 2006/05/06 01:56:44 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_clkgen_rtl_c0 of t400_clkgen is

  for rtl
  end for;

end t400_clkgen_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_clkgen-c.vhd,v $
-- Revision 1.1.1.1  2006/05/06 01:56:44  arniml
-- import from local CVS repository, LOC_CVS_0_1
--
-------------------------------------------------------------------------------
