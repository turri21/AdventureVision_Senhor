-------------------------------------------------------------------------------
--
-- The Data memory controller.
--
-- $Id: t400_dmem_ctrl-c.vhd,v 1.1.1.1 2006/05/06 01:56:44 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_dmem_ctrl_rtl_c0 of t400_dmem_ctrl is

  for rtl
  end for;

end t400_dmem_ctrl_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_dmem_ctrl-c.vhd,v $
-- Revision 1.1.1.1  2006/05/06 01:56:44  arniml
-- import from local CVS repository, LOC_CVS_0_1
--
-------------------------------------------------------------------------------
