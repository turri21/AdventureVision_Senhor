-------------------------------------------------------------------------------
--
-- The opcode decoder table.
-- Maps the binary opcodes to the mnemonic type.
--
-- $Id: t400_opc_table-c.vhd,v 1.1.1.1 2006/05/06 01:56:44 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_opc_table_rtl_c0 of t400_opc_table is

  for rtl
  end for;

end t400_opc_table_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: t400_opc_table-c.vhd,v $
-- Revision 1.1.1.1  2006/05/06 01:56:44  arniml
-- import from local CVS repository, LOC_CVS_0_1
--
-------------------------------------------------------------------------------
